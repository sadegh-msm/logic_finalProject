/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2021-2022
--  *******************************************************
--  Student ID  : 
--  Student Name: 
--  Student Mail: 
--  *******************************************************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: calculate_new_capacity
-----------------------------------------------------------*/
`timescale 1 ns/1 ns

module calculate_new_capacity(
	park_location,
	parking_capacity,
	new_capacity);
	
	input [7:0] park_location;
	input [7:0] parking_capacity;
	output reg [7:0] new_capacity;

	always @ (parking_capacity or park_location)
	begin
		new_capacity = park_location ^ parking_capacity;
	end
	
endmodule